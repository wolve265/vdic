interface alu_bfm;
	import alu_pkg::*;
	
	bit clk;
	bit rst_n;
	bit sin;
	bit sout;
	
endinterface : alu_bfm