module coverage(alu_bfm bfm);
	import alu_pkg::*;
	
endmodule : coverage