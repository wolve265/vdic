module tester(alu_bfm bfm);
	import alu_pkg::*;
	
endmodule : tester