package alu_pkg;
	
endpackage : alu_pkg