module scoreboard(alu_bfm bfm);
	import alu_pkg::*;
	
endmodule : scoreboard