
module top;
	
	initial begin : top_core
		$display("test");
	end : top_core
	
endmodule : top